
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity lfsr_testbench is
end lfsr_testbench;

architecture tb of lfsr_testbench is

	function vec2str(vec: std_logic_vector) return string is
    variable stmp: string(vec'left+1 downto 1);
    begin
        for i in vec'reverse_range loop
            if (vec(i) = 'U') then
                stmp(i+1) := 'U';
            elsif (vec(i) = 'X') then
                stmp(i+1) := 'X';
            elsif (vec(i) = '0') then
                stmp(i+1) := '0';
            elsif (vec(i) = '1') then
                stmp(i+1) := '1';
            elsif (vec(i) = 'Z') then
                stmp(i+1) := 'Z';
            elsif (vec(i) = 'W') then
                stmp(i+1) := 'W';
            elsif (vec(i) = 'L') then
                stmp(i+1) := 'L';
           elsif (vec(i) = 'H') then
                stmp(i+1) := 'H';
            else
                stmp(i+1) := '-';
            end if;
        end loop;
    return stmp;
    end;
	
	component lfsr
        generic (N    : integer;
                 SEED : std_logic_vector(130 downto 0));
        port (clk   : in std_logic;
              reset : in std_logic;
              q     : out std_logic_vector(130 downto 0));
    end component;

	signal lfsr_out1,lfsr_out2: std_logic_vector(130 downto 0);
	signal clk,rst: std_logic;

	constant period_t: time:=10 ns;
	constant period: integer:=10;
	--patterns generated by the lfsr's
	constant patterns: integer:=1000;
	--cycles needed
	constant cycles: integer:=patterns*(2*period);
    
begin

	uut_lfsr1: lfsr
	generic map(
		N=>130,
		SEED=>std_logic_vector(to_unsigned(1,131))
	)
	port map(
		clk=>clk,
		reset=>rst,
		q=>lfsr_out1
	);

	uut_lfsr2: lfsr
	generic map(
		N=>130,
		SEED=>std_logic_vector(to_unsigned(2,131))
	)
	port map(
		clk=>clk,
		reset=>rst,
		q=>lfsr_out2
	);
	

	process
	begin
		clk<='0';
		wait for period_t;
		clk<='1';
		wait for period_t;
	end process;

	process
	begin
		rst<='1';
		wait for 2 ns;
		rst<='0';
		wait;
	end process;

	process(clk)
	type patterns_array is array(0 to patterns-1) of std_logic_vector(130 downto 0);
	variable patterns1: patterns_array;
	variable patterns2: patterns_array;
	variable cycle_count: integer:=0;
	variable match_counter: integer :=0;
	variable i,j: integer:=0;
	begin
		if cycle_count=(patterns-1) then
			--compare
			for i in 0 to patterns-1 loop
				for j in 0 to patterns-1 loop 
					if patterns1(i) = patterns2(j) then
						match_counter:=match_counter+1;
						report "i "& integer'image(i) & " j " & integer'image(j);
						report "Pattern 1 "& vec2str(patterns1(i)) & " Is equal to pattern 2 " & vec2str(patterns2(j)) & CR & LF;
					end if;
				end loop;
			end loop;
			cycle_count:=patterns;
			assert false report "Found matches "& integer'image(match_counter) severity warning;
		elsif cycle_count < (patterns-1) then
			if rising_edge(clk) then
				patterns1(cycle_count):=lfsr_out1;
				patterns2(cycle_count):=lfsr_out2;
				cycle_count:=cycle_count + 1;
			end if;
		end if;
		
	end process;

end tb;

configuration cfg_lfsr_testbench of lfsr_testbench is
    for tb
    end for;
end cfg_lfsr_testbench;
