package constants is
    constant N_MISR: integer := 64;
end package constants;