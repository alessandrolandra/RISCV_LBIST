package constants is
    constant N_MISR: integer := 64;
	constant PATT_PATH_LOAD: string:= "./atpg_pat_converter/t_patterns.txt";
	constant PATT_PATH_CAP: string:= "./atpg_pat_converter/c_patterns.txt";
end package constants;
